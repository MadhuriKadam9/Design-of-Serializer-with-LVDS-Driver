* D:\Serializer_Lvds_dvr\PISO\PISO.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/10/22 16:00:41

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_U5-Pad5_ Net-_U5-Pad6_ Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_U5-Pad9_ Net-_U5-Pad10_ Net-_U5-Pad11_ Net-_U5-Pad12_ Net-_U10-Pad1_ madhuri_piso		
U8  clk load I9 GND I7 GND Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_U5-Pad5_ Net-_U5-Pad6_ adc_bridge_6		
U9  I5 GND I3 I2 I1 I0 Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_U5-Pad9_ Net-_U5-Pad10_ Net-_U5-Pad11_ Net-_U5-Pad12_ adc_bridge_6		
v1  clk GND pulse		
v2  load GND pulse		
v3  I3 GND pulse		
v4  I2 GND pulse		
v5  I1 GND pulse		
v6  I0 GND pulse		
U1  clk plot_v1		
U4  load plot_v1		
U3  I3 plot_v1		
U6  I2 plot_v1		
U2  I1 plot_v1		
U7  I0 plot_v1		
U11  Din plot_v1		
v9  I5 GND pulse		
v8  I7 GND pulse		
v7  I9 GND pulse		
U12  I9 plot_v1		
U13  I7 plot_v1		
U14  I5 plot_v1		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ madhuri_buffer		
U15  Din_bar plot_v1		
U16  Net-_U10-Pad2_ Net-_U10-Pad3_ Din Din_bar dac_bridge_2		

.end
